`timescale 10ns / 1ns
`include "interfaces.svh"

module test_app (
);

endmodule