`timescale 10ns / 1ns
`include "interfaces.svh"

module test_app_tb ();


endmodule